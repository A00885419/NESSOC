/*
	apu.sv
	audio processing unit
	This thing is a stretch goal but here is the dummy module anyway
*/

module apu(
	input logic [7:0] P1CTL,
	input logic [7:0] P1RAMP,
	input logic [7:0] P1FT,
	input logic [7:0] P1CT,
	input logic [7:0] P2CTL,
	input logic [7:0] P2RAMP,
	input logic [7:0] P2FT,
	input logic [7:0] P2FT,
	
);

endmodule