/*
vga.sv 

This is the vga output module

By writing to the frame buffer, the vga output is updated.

frame buffer -> vga out
*/

module vga(input );